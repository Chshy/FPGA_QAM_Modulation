module top (
    input clk,
    input rst_n
    // ports
);



    
endmodule
