module calc_step (
    input  [15:0] freq,
    output [ 9:0] step
);

// clk = 11.05926 MHz / 4
// f_sine = f_clk * 2^W / step
// step = f_clk * 4096 / f_sine

assign step = 
    freq < 16'd  507 ? 10'd   1 : 
    freq < 16'd  845 ? 10'd   2 : 
    freq < 16'd 1183 ? 10'd   3 : 
    freq < 16'd 1521 ? 10'd   4 : 
    freq < 16'd 1859 ? 10'd   5 : 
    freq < 16'd 2197 ? 10'd   6 : 
    freq < 16'd 2535 ? 10'd   7 : 
    freq < 16'd 2873 ? 10'd   8 : 
    freq < 16'd 3211 ? 10'd   9 : 
    freq < 16'd 3549 ? 10'd  10 : 
    freq < 16'd 3887 ? 10'd  11 : 
    freq < 16'd 4225 ? 10'd  12 : 
    freq < 16'd 4563 ? 10'd  13 : 
    freq < 16'd 4901 ? 10'd  14 : 
    freq < 16'd 5239 ? 10'd  15 : 
    freq < 16'd 5577 ? 10'd  16 : 
    freq < 16'd 5915 ? 10'd  17 : 
    freq < 16'd 6253 ? 10'd  18 : 
    freq < 16'd 6591 ? 10'd  19 : 
    freq < 16'd 6929 ? 10'd  20 : 
    freq < 16'd 7267 ? 10'd  21 : 
    freq < 16'd 7605 ? 10'd  22 : 
    freq < 16'd 7943 ? 10'd  23 : 
    freq < 16'd 8281 ? 10'd  24 : 
    freq < 16'd 8619 ? 10'd  25 : 
    freq < 16'd 8957 ? 10'd  26 : 
    freq < 16'd 9295 ? 10'd  27 : 
    freq < 16'd 9633 ? 10'd  28 : 
    freq < 16'd 9971 ? 10'd  29 : 
    freq < 16'd10309 ? 10'd  30 : 
    freq < 16'd10647 ? 10'd  31 : 
    freq < 16'd10985 ? 10'd  32 : 
    freq < 16'd11323 ? 10'd  33 : 
    freq < 16'd11661 ? 10'd  34 : 
    freq < 16'd11999 ? 10'd  35 : 
    freq < 16'd12337 ? 10'd  36 : 
    freq < 16'd12675 ? 10'd  37 : 
    freq < 16'd13013 ? 10'd  38 : 
    freq < 16'd13351 ? 10'd  39 : 
    freq < 16'd13689 ? 10'd  40 : 
    freq < 16'd14027 ? 10'd  41 : 
    freq < 16'd14365 ? 10'd  42 : 
    freq < 16'd14703 ? 10'd  43 : 
    freq < 16'd15041 ? 10'd  44 : 
    freq < 16'd15379 ? 10'd  45 : 
    freq < 16'd15717 ? 10'd  46 : 
    freq < 16'd16055 ? 10'd  47 : 
    freq < 16'd16393 ? 10'd  48 : 
    freq < 16'd16731 ? 10'd  49 : 
    freq < 16'd17069 ? 10'd  50 : 
    freq < 16'd17407 ? 10'd  51 : 
    freq < 16'd17745 ? 10'd  52 : 
    freq < 16'd18083 ? 10'd  53 : 
    freq < 16'd18421 ? 10'd  54 : 
    freq < 16'd18759 ? 10'd  55 : 
    freq < 16'd19097 ? 10'd  56 : 
    freq < 16'd19435 ? 10'd  57 : 
    freq < 16'd19773 ? 10'd  58 : 
    freq < 16'd20111 ? 10'd  59 : 
    freq < 16'd20449 ? 10'd  60 : 
    freq < 16'd20787 ? 10'd  61 : 
    freq < 16'd21125 ? 10'd  62 : 
    freq < 16'd21463 ? 10'd  63 : 
    freq < 16'd21801 ? 10'd  64 : 
    freq < 16'd22139 ? 10'd  65 : 
    freq < 16'd22477 ? 10'd  66 : 
    freq < 16'd22815 ? 10'd  67 : 
    freq < 16'd23153 ? 10'd  68 : 
    freq < 16'd23491 ? 10'd  69 : 
    freq < 16'd23829 ? 10'd  70 : 
    freq < 16'd24167 ? 10'd  71 : 
    freq < 16'd24505 ? 10'd  72 : 
    freq < 16'd24843 ? 10'd  73 : 
    freq < 16'd25181 ? 10'd  74 : 
    freq < 16'd25519 ? 10'd  75 : 
    freq < 16'd25857 ? 10'd  76 : 
    freq < 16'd26195 ? 10'd  77 : 
    freq < 16'd26533 ? 10'd  78 : 
    freq < 16'd26871 ? 10'd  79 : 
    freq < 16'd27209 ? 10'd  80 : 
    freq < 16'd27547 ? 10'd  81 : 
    freq < 16'd27885 ? 10'd  82 : 
    freq < 16'd28223 ? 10'd  83 : 
    freq < 16'd28561 ? 10'd  84 : 
    freq < 16'd28899 ? 10'd  85 : 
    freq < 16'd29237 ? 10'd  86 : 
    freq < 16'd29575 ? 10'd  87 : 
    freq < 16'd29913 ? 10'd  88 : 
    freq < 16'd30251 ? 10'd  89 : 
    freq < 16'd30589 ? 10'd  90 : 
    freq < 16'd30927 ? 10'd  91 : 
    freq < 16'd31265 ? 10'd  92 : 
    freq < 16'd31603 ? 10'd  93 : 
    freq < 16'd31941 ? 10'd  94 : 
    freq < 16'd32279 ? 10'd  95 : 
    freq < 16'd32617 ? 10'd  96 : 
    freq < 16'd32955 ? 10'd  97 : 
    freq < 16'd33293 ? 10'd  98 : 
    freq < 16'd33631 ? 10'd  99 : 
    freq < 16'd33969 ? 10'd 100 : 
    freq < 16'd34307 ? 10'd 101 : 
    freq < 16'd34645 ? 10'd 102 : 
    freq < 16'd34983 ? 10'd 103 : 
    freq < 16'd35321 ? 10'd 104 : 
    freq < 16'd35659 ? 10'd 105 : 
    freq < 16'd35997 ? 10'd 106 : 
    freq < 16'd36335 ? 10'd 107 : 
    freq < 16'd36673 ? 10'd 108 : 
    freq < 16'd37011 ? 10'd 109 : 
    freq < 16'd37349 ? 10'd 110 : 
    freq < 16'd37687 ? 10'd 111 : 
    freq < 16'd38025 ? 10'd 112 : 
    freq < 16'd38363 ? 10'd 113 : 
    freq < 16'd38701 ? 10'd 114 : 
    freq < 16'd39039 ? 10'd 115 : 
    freq < 16'd39377 ? 10'd 116 : 
    freq < 16'd39715 ? 10'd 117 : 
    freq < 16'd40053 ? 10'd 118 : 
    freq < 16'd40391 ? 10'd 119 : 
    freq < 16'd40729 ? 10'd 120 : 
    freq < 16'd41067 ? 10'd 121 : 
    freq < 16'd41405 ? 10'd 122 : 
    freq < 16'd41743 ? 10'd 123 : 
    freq < 16'd42081 ? 10'd 124 : 
    freq < 16'd42419 ? 10'd 125 : 
    freq < 16'd42757 ? 10'd 126 : 
    freq < 16'd43095 ? 10'd 127 : 
    freq < 16'd43433 ? 10'd 128 : 
    freq < 16'd43771 ? 10'd 129 : 
    freq < 16'd44109 ? 10'd 130 : 
    freq < 16'd44447 ? 10'd 131 : 
    freq < 16'd44785 ? 10'd 132 : 
    freq < 16'd45123 ? 10'd 133 : 
    freq < 16'd45461 ? 10'd 134 : 
    freq < 16'd45799 ? 10'd 135 : 
    freq < 16'd46137 ? 10'd 136 : 
    freq < 16'd46475 ? 10'd 137 : 
    freq < 16'd46813 ? 10'd 138 : 
    freq < 16'd47151 ? 10'd 139 : 
    freq < 16'd47489 ? 10'd 140 : 
    freq < 16'd47827 ? 10'd 141 : 
    freq < 16'd48165 ? 10'd 142 : 
    freq < 16'd48503 ? 10'd 143 : 
    freq < 16'd48841 ? 10'd 144 : 
    freq < 16'd49179 ? 10'd 145 : 
    freq < 16'd49517 ? 10'd 146 : 
    freq < 16'd49855 ? 10'd 147 : 
    freq < 16'd50193 ? 10'd 148 : 
    freq < 16'd50531 ? 10'd 149 : 
    freq < 16'd50869 ? 10'd 150 : 
    freq < 16'd51207 ? 10'd 151 : 
    freq < 16'd51545 ? 10'd 152 : 
    freq < 16'd51883 ? 10'd 153 : 
    freq < 16'd52221 ? 10'd 154 : 
    freq < 16'd52559 ? 10'd 155 : 
    freq < 16'd52897 ? 10'd 156 : 
    freq < 16'd53235 ? 10'd 157 : 
    freq < 16'd53573 ? 10'd 158 : 
    freq < 16'd53911 ? 10'd 159 : 
    freq < 16'd54249 ? 10'd 160 : 
    freq < 16'd54587 ? 10'd 161 : 
    freq < 16'd54925 ? 10'd 162 : 
    freq < 16'd55263 ? 10'd 163 : 
    freq < 16'd55601 ? 10'd 164 : 
    freq < 16'd55939 ? 10'd 165 : 
    freq < 16'd56277 ? 10'd 166 : 
    freq < 16'd56615 ? 10'd 167 : 
    freq < 16'd56953 ? 10'd 168 : 
    freq < 16'd57291 ? 10'd 169 : 
    freq < 16'd57629 ? 10'd 170 : 
    freq < 16'd57967 ? 10'd 171 : 
    freq < 16'd58305 ? 10'd 172 : 
    freq < 16'd58643 ? 10'd 173 : 
    freq < 16'd58981 ? 10'd 174 : 
    freq < 16'd59319 ? 10'd 175 : 
    freq < 16'd59657 ? 10'd 176 : 
    freq < 16'd59995 ? 10'd 177 : 
    freq < 16'd60333 ? 10'd 178 : 
    freq < 16'd60671 ? 10'd 179 : 
    freq < 16'd61009 ? 10'd 180 : 
    freq < 16'd61347 ? 10'd 181 : 
    freq < 16'd61685 ? 10'd 182 : 
    freq < 16'd62023 ? 10'd 183 : 
    freq < 16'd62361 ? 10'd 184 : 
    freq < 16'd62699 ? 10'd 185 : 
    freq < 16'd63037 ? 10'd 186 : 
    freq < 16'd63375 ? 10'd 187 : 
    freq < 16'd63713 ? 10'd 188 : 
    freq < 16'd64051 ? 10'd 189 : 
    freq < 16'd64389 ? 10'd 190 : 
    freq < 16'd64727 ? 10'd 191 : 
    freq < 16'd65065 ? 10'd 192 : 
    freq < 16'd65403 ? 10'd 193 : 
                       10'd 194 ;
endmodule